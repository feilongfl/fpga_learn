/////////////////////////////////////////////
// author: feilong
// version: 1.0.0
/////////////////////////////////////////////

module divclk (
           input  clk_in,
           output reg clk_out
       );
/////////////////////////////////////////////
// parameter and signals
/////////////////////////////////////////////
// parameter
parameter DIV_COUNT = 10;

// regs or wires
reg[15:0] count = 0;
/////////////////////////////////////////////
// main code
/////////////////////////////////////////////

always @ (posedge clk_in) begin
    count <= (count == DIV_COUNT - 1)? 0 : count + 1;
end

always @ (posedge clk_in) begin
    clk_out <= (count < (DIV_COUNT / 2)) ? 1 : 0;
end

/////////////////////////////////////////////
// code end
/////////////////////////////////////////////
endmodule
