/////////////////////////////////////////////
// author: feilong
// version: 1.0.0
/////////////////////////////////////////////

module recviver (
           input  clk,
           input  en,
           input  rx,
           output reg [7:0]data
       );
/////////////////////////////////////////////
// parameter and signals
/////////////////////////////////////////////
// parameter

// regs or wires

/////////////////////////////////////////////
// main code
/////////////////////////////////////////////



/////////////////////////////////////////////
// code end
/////////////////////////////////////////////
endmodule
