/////////////////////////////////////////////
// author: feilong
// version: 1.0.0
/////////////////////////////////////////////

module ddrAddrGen (
           input  flags,
           output reg [27:0] Addr = 0,
           output reg [31:0] mask = 32'b11111111_11111111_11111111_11111110
       );
/////////////////////////////////////////////
// parameter and signals
/////////////////////////////////////////////
// parameter

// regs or wires

/////////////////////////////////////////////
// main code
/////////////////////////////////////////////
always @ (posedge flags) begin
    mask <= (mask == 32'b01111111_11111111_11111111_11111111)?
         32'b11111111_11111111_11111111_11111110 : (mask << 1);

    Addr <= (mask == 32'b01111111_11111111_11111111_11111111)? Addr + 1 : Addr;
end


/////////////////////////////////////////////
// code end
/////////////////////////////////////////////
endmodule
