/////////////////////////////////////////////
// author: feilong
// version: 1.0.0
/////////////////////////////////////////////

module signalChangeDector (
           input  clk,
           input signal,
           output trig
       );
/////////////////////////////////////////////
// parameter and signals
/////////////////////////////////////////////
// parameter
parameter BufferSize = 2;
parameter BufferInital = 0;
// regs or wires
reg [BufferSize : 0] buff = BufferInital;
/////////////////////////////////////////////
// main code
/////////////////////////////////////////////
always @ (posedge clk) begin
    buff <= {buff[BufferSize - 1 : 0],signal};
end

assign trig = (buff[BufferSize] == buff[BufferSize - 1])? 0 : 1;
/////////////////////////////////////////////
// code end
/////////////////////////////////////////////
endmodule
