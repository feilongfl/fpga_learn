/////////////////////////////////////////////
// author: feilong
// version: 1.0.0
/////////////////////////////////////////////

module writeRamAddrGen (
           input enable,
           input  rxflag,

           input[7:0] dataLength,

           output reg [7:0] ramAddress = 0,
           output reg finishFlag = 0
       );
/////////////////////////////////////////////
// parameter and signals
/////////////////////////////////////////////
// parameter

// regs or wires

/////////////////////////////////////////////
// main code
/////////////////////////////////////////////
always @ (posedge rxflag) begin
    ramAddress <= (enable)? ramAddress + 1 : 0;

    finishFlag <= (ramAddress + 1 == dataLength)? 1 : 0;
end

/////////////////////////////////////////////
// code end
/////////////////////////////////////////////
endmodule
