/////////////////////////////////////////////
// author: feilong
// version: 1.0.0
/////////////////////////////////////////////

module bit8mask256 (
           input [7:0] I,
           // input [31:0]mask,
           output [255:0] O
       );
/////////////////////////////////////////////
// parameter and signals
/////////////////////////////////////////////
// parameter

// regs or wires
// wire[31:0] notMask;

/////////////////////////////////////////////
// main code
/////////////////////////////////////////////
// assign notMask = ~(mask);
assign O = {
           I,I,I,I,I,I,I,I,
           I,I,I,I,I,I,I,I,
           I,I,I,I,I,I,I,I,
           I,I,I,I,I,I,I,I
       };


/////////////////////////////////////////////
// code end
/////////////////////////////////////////////
endmodule
