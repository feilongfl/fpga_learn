/////////////////////////////////////////////
// author: feilong
// version: 1.0.0
/////////////////////////////////////////////

module recv_clk_gen (
           input  rx,
           input clk,
           output outval
       );
/////////////////////////////////////////////
// parameter and signals
/////////////////////////////////////////////
// parameter
parameter TIME_MAX = 5206;
parameter TRIG_AT = TIME_MAX / 2;
parameter TRIG_TIME = 10;

// regs or wires
reg[31:0] count = 0;
reg en = 0;
/////////////////////////////////////////////
// main code
/////////////////////////////////////////////
always @ (negedge rx) begin
    en = 1;
end


always @ (posedge clk) begin
    count <= (count == TIME_MAX)? 0 : count + 1;
end


/////////////////////////////////////////////
// code end
/////////////////////////////////////////////
endmodule
