/////////////////////////////////////////////
// author: feilong
// version: 1.0.0
/////////////////////////////////////////////

module fifo (
           input  clk,
           input  indata,
           output outdata
       );
/////////////////////////////////////////////
// parameter and signals
/////////////////////////////////////////////
// parameter

// regs or wires
reg[2:0] data_buff = 0;
/////////////////////////////////////////////
// main code
/////////////////////////////////////////////
always @ (posedge clk) begin
    data_buff <= {data_buff[1:0],indata};
end

assign outdata = data_buff[2];

/////////////////////////////////////////////
// code end
/////////////////////////////////////////////
endmodule
