/////////////////////////////////////////////
// author: feilong
// version: 1.0.0
/////////////////////////////////////////////

module top (
	    input 	 clk,
	    input 	 rst,
	    input 	 button,
	    output [3:0] leds
	    );
	/////////////////////////////////////////////
	// parameter and signals
	/////////////////////////////////////////////
	// parameter

	// regs or wires
	wire 		 button_sig;
	/////////////////////////////////////////////
	// main code
	/////////////////////////////////////////////
	led led_inst(
    		     .iclk(button_sig),
    		     .rst(rst),
    		     .leds(leds)
    		     );

	button button_inst(
			   .clk(clk),
			   .button_in(button),
			   .button_out(button_sig)
			   );


	/////////////////////////////////////////////
	// code end
	/////////////////////////////////////////////
endmodule
