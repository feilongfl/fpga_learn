/////////////////////////////////////////////
// author: feilong
// version: 1.0.0
/////////////////////////////////////////////

module modulename (
		   input  inval,
		   output outval
		   );
    /////////////////////////////////////////////
    // parameter and signals
    /////////////////////////////////////////////
    // parameter

    // regs

    /////////////////////////////////////////////
    // main code
    /////////////////////////////////////////////



    /////////////////////////////////////////////
    // code end
    /////////////////////////////////////////////
endmodule
