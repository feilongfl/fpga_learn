/////////////////////////////////////////////
// author: feilong
// version: 1.0.0
/////////////////////////////////////////////

module top (
           input  sclk,
           input srst_r,
           output hsync,vsync,
           output r,g,b
       );
/////////////////////////////////////////////
// parameter and signals
/////////////////////////////////////////////
// parameter

// regs or wires

/////////////////////////////////////////////
// main code
/////////////////////////////////////////////



/////////////////////////////////////////////
// code end
/////////////////////////////////////////////
endmodule
