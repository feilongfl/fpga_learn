/////////////////////////////////////////////
// author: feilong
// version: 1.0.0
/////////////////////////////////////////////

module uart (
           input  uart_rx,
           output uart_tx,

           // input[7:0] data_send,
           // input data_send_trig,
           output[7:0] data_recv,
           output data_recv_flag,

           input clock
       );
/////////////////////////////////////////////
// parameter and signals
/////////////////////////////////////////////
// parameter
parameter bandRate = 115200;
parameter clockSpeed = 50_000_000;
// regs or wires

/////////////////////////////////////////////
// main code
/////////////////////////////////////////////



/////////////////////////////////////////////
// code end
/////////////////////////////////////////////
endmodule
