/////////////////////////////////////////////
// author: feilong
// version: 1.0.0
/////////////////////////////////////////////

module cov1_8 (
           input  i,
           output [7:0] o
       );
/////////////////////////////////////////////
// parameter and signals
/////////////////////////////////////////////
// parameter

// regs or wires

/////////////////////////////////////////////
// main code
/////////////////////////////////////////////
assign o = {i,i,i,i,i,i,i,i};



/////////////////////////////////////////////
// code end
/////////////////////////////////////////////
endmodule
