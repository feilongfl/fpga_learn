
module vio (
	source);	

	output	[0:0]	source;
endmodule
