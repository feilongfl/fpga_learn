/////////////////////////////////////////////
// author: feilong
// version: 1.0.0
/////////////////////////////////////////////

module datasaver (
           input  saveflag,
           input [7:0]data_i,
           output reg [7:0] data_o = 0
       );
/////////////////////////////////////////////
// parameter and signals
/////////////////////////////////////////////
// parameter

// regs or wires

/////////////////////////////////////////////
// main code
/////////////////////////////////////////////

always @ (posedge saveflag) begin
    data_o <= data_i;
end

/////////////////////////////////////////////
// code end
/////////////////////////////////////////////
endmodule
