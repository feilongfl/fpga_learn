/////////////////////////////////////////////
// author: feilong
// version: 1.0.0
/////////////////////////////////////////////

module ddrctl (
           input  inval,
           output outval
       );
/////////////////////////////////////////////
// parameter and signals
/////////////////////////////////////////////
// parameter

// regs or wires

/////////////////////////////////////////////
// main code
/////////////////////////////////////////////



/////////////////////////////////////////////
// code end
/////////////////////////////////////////////
endmodule
