/////////////////////////////////////////////
// author: feilong
// version: 1.0.0
/////////////////////////////////////////////

module drinkouter (
		   input  en,
		   output drink_contral
		   );
	/////////////////////////////////////////////
	// parameter and signals
	/////////////////////////////////////////////
	// parameter

	// regs or wires

	/////////////////////////////////////////////
	// main code
	/////////////////////////////////////////////
	assign drink_contral = en;

	/////////////////////////////////////////////
	// code end
	/////////////////////////////////////////////
endmodule
