/////////////////////////////////////////////
// author: feilong
// version: 1.0.0
/////////////////////////////////////////////

module color (
           input  [15:0]x,
           input  [15:0]y,
           output [7:0]r,
           output [7:0]g,
           output [7:0]b
       );
/////////////////////////////////////////////
// parameter and signals
/////////////////////////////////////////////
// parameter
parameter eage1 = 160;
parameter eage2 = 320;

// regs or wires

/////////////////////////////////////////////
// main code
/////////////////////////////////////////////
assign r = (y < eage1) ? 8'hff : 0;
assign g = (y < eage2 && y >= eage1) ? 8'hff : 0;
assign b = (y >= eage2) ? 8'hff : 0;



/////////////////////////////////////////////
// code end
/////////////////////////////////////////////
endmodule
