/////////////////////////////////////////////
// author: feilong
// version: 1.0.0
/////////////////////////////////////////////

module SignalDelay (
           input  clk,
           input signal,
           output signalOut
       );
/////////////////////////////////////////////
// parameter and signals
/////////////////////////////////////////////
// parameter
parameter length = 1;
// regs or wires
reg [length:0] Buff = 0;
/////////////////////////////////////////////
// main code
/////////////////////////////////////////////
always @ (posedge clk) begin
    Buff <= {Buff[length - 1 : 0],signal};
end

assign signalOut = Buff[length];
/////////////////////////////////////////////
// code end
/////////////////////////////////////////////
endmodule
