/////////////////////////////////////////////
// author: feilong
// version: 1.0.0
/////////////////////////////////////////////

module cov8_1 (
           input [7:0] i,
           output o
       );
/////////////////////////////////////////////
// parameter and signals
/////////////////////////////////////////////
// parameter

// regs or wires

/////////////////////////////////////////////
// main code
/////////////////////////////////////////////
assign o = i[0] | i[1] | i[2] | i[3] | i[4] | i[5] | i[6] | i[7];



/////////////////////////////////////////////
// code end
/////////////////////////////////////////////
endmodule
