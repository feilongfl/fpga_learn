/////////////////////////////////////////////
// author: feilong
// version: 1.0.0
/////////////////////////////////////////////

module white (
           output r,g,b
       );
/////////////////////////////////////////////
// parameter and signals
/////////////////////////////////////////////
// parameter

// regs or wires

/////////////////////////////////////////////
// main code
/////////////////////////////////////////////
assign r = 1'b1;
assign g = 1'b1;
assign b = 1'b1;

/////////////////////////////////////////////
// code end
/////////////////////////////////////////////
endmodule
