/////////////////////////////////////////////
// author: feilong
// version: 1.0.0
/////////////////////////////////////////////

module color_flash (
           input clk,
           input [7:0] data,
           output [7:0] r,g,b
       );
/////////////////////////////////////////////
// parameter and signals
/////////////////////////////////////////////
// parameter

// regs or wires
reg [2:0] cnt = 0;
/////////////////////////////////////////////
// main code
/////////////////////////////////////////////
always @ (posedge clk) begin
    cnt <= (cnt == 5)? 0 : cnt + 1;
end

assign r = (cnt == 0 || cnt == 1 || cnt == 5)? data : 0;
assign g = (cnt == 1 || cnt == 2|| cnt == 3)? data : 0;
assign b = (cnt == 3 || cnt == 4 || cnt == 5)? data : 0;


/////////////////////////////////////////////
// code end
/////////////////////////////////////////////
endmodule
