/////////////////////////////////////////////
// author: feilong
// version: 1.0.0
/////////////////////////////////////////////

module led (
	    input 	     iclk,
	    input 	     rst,
	    output reg [3:0] leds
	    );
	/////////////////////////////////////////////
	// parameter and signals
	/////////////////////////////////////////////
	// parameter

	// regs

	/////////////////////////////////////////////
	// main code
	/////////////////////////////////////////////
	always @ (posedge iclk or negedge rst) begin
		if (!rst) begin
			leds <= 4'b0001;
		end else begin
			leds <= {leds[2:0],leds[3]};
		end
	end


	/////////////////////////////////////////////
	// code end
	/////////////////////////////////////////////
endmodule
