/////////////////////////////////////////////
// author: feilong
// version: 1.0.0
/////////////////////////////////////////////

module drinkouter (
		   input      en,
		   input      drink_out_fin,
		   output     drink_contral,
		   output reg flag = 1
		   );
	/////////////////////////////////////////////
	// parameter and signals
	/////////////////////////////////////////////
	// parameter

	// regs or wires

	/////////////////////////////////////////////
	// main code
	/////////////////////////////////////////////
	assign drink_contral = ~(en & flag);
	always @ (posedge en or negedge drink_out_fin) begin
		if(!drink_out_fin)
			flag <= 0;
		else
			flag <= 1;
	end
	/////////////////////////////////////////////
	// code end
	/////////////////////////////////////////////
endmodule
