typedef enum bit [4:0] {
	S_SDRAM_Initial,
	S_SDRAM_ARBIT,
	S_SDRAM_AutoRefresh,
	S_SDRAM_Write_once,
	S_SDRAM_READ
} StatusSdram_t;
