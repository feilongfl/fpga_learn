/////////////////////////////////////////////
// author: feilong
// version: 1.0.0
/////////////////////////////////////////////

module divclk (
           input  iclk,
           output oclk
       );
/////////////////////////////////////////////
// parameter and signals
/////////////////////////////////////////////
// parameter
parameter DIV_COUNT_MAX = 9;

// regs or wires
reg[4:0] count = 0;
/////////////////////////////////////////////
// main code
/////////////////////////////////////////////
always @ (posedge iclk) begin
    count <= count + 1;
end

assign oclk = (count < (DIV_COUNT_MAX + 1) / 2) ? 1 : 0;


/////////////////////////////////////////////
// code end
/////////////////////////////////////////////
endmodule
