/////////////////////////////////////////////
// author: feilong
// version: 1.0.0
/////////////////////////////////////////////

module pos_neg_dector (
           input  insig,
           input clk,
           output trig
       );
/////////////////////////////////////////////
// parameter and signals
/////////////////////////////////////////////
// parameter
parameter initial_val = 0;
// regs or wires
reg insig_last = initial_val;
/////////////////////////////////////////////
// main code
/////////////////////////////////////////////
always @ (posedge clk) begin
    insig_last <= insig;
end

assign trig = insig ^ insig_last;
/////////////////////////////////////////////
// code end
/////////////////////////////////////////////
endmodule
